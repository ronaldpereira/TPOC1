`include "alu.v"

module testbench;

	reg clock = 0, clear = 0;
	reg [31:0] inputA, inputB;
	reg [2:0] opCode;
	wire zero;
	wire [31:0] result;

	always #1 clock = !clock;

	initial $dumpfile("testbench.vcd");
	initial $dumpvars(0, testbench);

	alu c(clock, clear, result, zero, inputA, inputB, opCode);

	initial
	begin
		#1 clear = 1;
		#1 clear = 0;
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000000100101110;
		#5 opCode = 3'b000; // 805 + 302 = 1107
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000000100101110;
		#5 opCode = 3'b001; // 805 - 302 = 503
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000001100100101;
		#5 opCode = 3'b001; // 805 - 805 = 0
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000001100100101;
		#5 opCode = 3'b010; // 805 AND 805 = 805
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000000100101110;
		#5 opCode = 3'b010; // 805 AND 302 = 292
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000000100101110;
		#5 opCode = 3'b011; // 805 OR 302 = 815
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000000100101110;
		#5 opCode = 3'b100; // 805 XOR 302 = 523
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000000100101110;
		#5 opCode = 3'b101; // 805 NOP 302 = 0
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000000100101110;
		#5 opCode = 3'b110; // 805 NOP 302 = 0
		#5 inputA = 32'b00000000000000000000001100100101;
		#5 inputB = 32'b00000000000000000000000100101110;
		#5 opCode = 3'b111; // 805 NOP 302 = 0
		#5 clear = 1;
		#5 $finish;
	end

endmodule // testbench
